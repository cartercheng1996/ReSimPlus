`timescale 1ns/1ps
module count(
   input        rst,
   input        clk,
   output [3:0] count_out);


endmodule
